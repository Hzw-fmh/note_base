module andd(
    input[3:0] A,B,
    output[3:0] res
);

assign res=A&B;
endmodule